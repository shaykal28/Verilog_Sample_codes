module clockbuffer(input in_clock,output buffered_clock);



buf one (buffered_clock,in_clock);

endmodule 